`default_nettype none

module top (
    input logic CLOCK_50, // 50 MHz
    input logic TD_RESET_N,

    output logic VGA_CLK,
    output logic [7:0] VGA_R,
    output logic [7:0] VGA_G,
    output logic [7:0] VGA_B,

    output logic VGA_SYNC_N, // sync when 0
    output logic VGA_BLANK_N, // output data when 1

    output logic VGA_HS,
    output logic VGA_VS,
    );

    // PLL
    clk25 PLL (
        .clk(CLOCK_50),
        .n_rst(TD_RESET_N),
        .clk_25(VGA_CLK)
    );

    // VGA Controller
    logic video_on;
    logic [9:0] x_coordinate;
    logic [9:0] y_coordinate;
    vga_controller VGA_CNT (
        .clk_25(VGA_CLK),
        .n_rst(TD_RESET_N),
        .hsync(VGA_HS),
        .vsync(VGA_VS),
        .video_on(VGA_BLANK_N),
        .x_coordinate(x_coordinate),
        .y_coordinate(y_coordinate)
    );

    // Output
    logic [23:0] pixel_data;
    memory MEM (
        .pixel_x(x_coordinate),
        .pixel_y(y_coordinate),
        .pixel_data(pixel_data)
    );

    load_image MONITOR (
        .load_enable(video_on),
        .pixel_data(pixel_data),
        .red(VGA_R),
        .green(VGA_G),
        .blue(VGA_B)
    );
    
endmodule
